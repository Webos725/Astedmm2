<svg xmlns="http://www.w3.org/2000/svg" width="100" height="100" viewBox="0 0 100 100">
  <g stroke="black" stroke-width="3" fill="none">
    <!-- 上部：亠 -->
    <circle cx="50" cy="20" r="4" />
    <line x1="40" y1="30" x2="60" y2="30" />
    
    <!-- 中央：中心者 -->
    <line x1="50" y1="30" x2="50" y2="70" />
    
    <!-- 下部：糸の束感 -->
    <line x1="40" y1="60" x2="60" y2="60" />
    <line x1="45" y1="70" x2="55" y2="70" />
  </g>
</svg>
